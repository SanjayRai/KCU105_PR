module PR_module_A (
    input clk,
    output [15:0] data_out
);

endmodule
